// $Id: $
// File name:   cycle_counter.sv
// Created:     11/30/2014
// Author:      Sheik Dawood
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Cycle counter

module cycle_counter(
		     input wire clk,
		     input wire n_rst,
		     input wire 
		     );

   counter #(6) cycle(.clk(),

endmodule // cycle_counter

